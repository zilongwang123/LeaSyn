module ALU_3stage(
  input  [3:0]  io_fn,
  input  [31:0] io_in2,
  input  [31:0] io_in1,
  output [31:0] io_out,
  output [31:0] io_adder_out
);
  wire [31:0] _sum_T_2 = 32'h0 - io_in2; // @[alu.scala 50:40]
  wire [31:0] _sum_T_3 = io_fn[3] ? _sum_T_2 : io_in2; // @[alu.scala 50:25]
  wire [31:0] sum = io_in1 + _sum_T_3; // @[alu.scala 50:20]
  wire  _less_T_7 = io_fn[1] ? io_in2[31] : io_in1[31]; // @[alu.scala 54:18]
  wire  less = io_in1[31] == io_in2[31] ? sum[31] : _less_T_7; // @[alu.scala 53:19]
  wire [4:0] shamt = io_in2[4:0]; // @[alu.scala 58:21]
  wire  _shin_T_2 = io_fn == 4'h5 | io_fn == 4'hb; // @[alu.scala 60:37]
  wire [31:0] _GEN_0 = {{16'd0}, io_in1[31:16]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_6 = _GEN_0 & 32'hffff; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_8 = {io_in1[15:0], 16'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_10 = _shin_T_8 & 32'hffff0000; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_11 = _shin_T_6 | _shin_T_10; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_1 = {{8'd0}, _shin_T_11[31:8]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_16 = _GEN_1 & 32'hff00ff; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_18 = {_shin_T_11[23:0], 8'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_20 = _shin_T_18 & 32'hff00ff00; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_21 = _shin_T_16 | _shin_T_20; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_2 = {{4'd0}, _shin_T_21[31:4]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_26 = _GEN_2 & 32'hf0f0f0f; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_28 = {_shin_T_21[27:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_30 = _shin_T_28 & 32'hf0f0f0f0; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_31 = _shin_T_26 | _shin_T_30; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_3 = {{2'd0}, _shin_T_31[31:2]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_36 = _GEN_3 & 32'h33333333; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_38 = {_shin_T_31[29:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_40 = _shin_T_38 & 32'hcccccccc; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_41 = _shin_T_36 | _shin_T_40; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_4 = {{1'd0}, _shin_T_41[31:1]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_46 = _GEN_4 & 32'h55555555; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_48 = {_shin_T_41[30:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_50 = _shin_T_48 & 32'haaaaaaaa; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_51 = _shin_T_46 | _shin_T_50; // @[Bitwise.scala 105:39]
  wire [31:0] shin = io_fn == 4'h5 | io_fn == 4'hb ? io_in1 : _shin_T_51; // @[alu.scala 60:17]
  wire  _shout_r_T_2 = io_fn[3] & shin[31]; // @[alu.scala 61:35]
  wire [32:0] _shout_r_T_4 = {_shout_r_T_2,shin}; // @[alu.scala 61:60]
  wire [32:0] _shout_r_T_5 = $signed(_shout_r_T_4) >>> shamt; // @[alu.scala 61:63]
  wire [31:0] shout_r = _shout_r_T_5[31:0]; // @[alu.scala 61:72]
  wire [31:0] _GEN_5 = {{16'd0}, shout_r[31:16]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_3 = _GEN_5 & 32'hffff; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_5 = {shout_r[15:0], 16'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_7 = _shout_l_T_5 & 32'hffff0000; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_6 = {{8'd0}, _shout_l_T_8[31:8]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_13 = _GEN_6 & 32'hff00ff; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_15 = {_shout_l_T_8[23:0], 8'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_17 = _shout_l_T_15 & 32'hff00ff00; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_7 = {{4'd0}, _shout_l_T_18[31:4]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_23 = _GEN_7 & 32'hf0f0f0f; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_25 = {_shout_l_T_18[27:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_27 = _shout_l_T_25 & 32'hf0f0f0f0; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_8 = {{2'd0}, _shout_l_T_28[31:2]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_33 = _GEN_8 & 32'h33333333; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_35 = {_shout_l_T_28[29:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_37 = _shout_l_T_35 & 32'hcccccccc; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_9 = {{1'd0}, _shout_l_T_38[31:1]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_43 = _GEN_9 & 32'h55555555; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_45 = {_shout_l_T_38[30:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_47 = _shout_l_T_45 & 32'haaaaaaaa; // @[Bitwise.scala 105:80]
  wire [31:0] shout_l = _shout_l_T_43 | _shout_l_T_47; // @[Bitwise.scala 105:39]
  wire [31:0] _bitwise_logic_T_1 = io_in1 & io_in2; // @[alu.scala 65:35]
  wire [31:0] _bitwise_logic_T_3 = io_in1 | io_in2; // @[alu.scala 66:35]
  wire [31:0] _bitwise_logic_T_5 = io_in1 ^ io_in2; // @[alu.scala 67:35]
  wire [31:0] _bitwise_logic_T_6 = io_fn == 4'h4 ? _bitwise_logic_T_5 : io_in1; // @[alu.scala 67:8]
  wire [31:0] _bitwise_logic_T_7 = io_fn == 4'h6 ? _bitwise_logic_T_3 : _bitwise_logic_T_6; // @[alu.scala 66:8]
  wire [31:0] bitwise_logic = io_fn == 4'h7 ? _bitwise_logic_T_1 : _bitwise_logic_T_7; // @[alu.scala 65:8]
  wire [31:0] _out_xpr_length_T_10 = io_fn == 4'h1 ? shout_l : bitwise_logic; // @[alu.scala 74:8]
  wire [31:0] _out_xpr_length_T_11 = _shin_T_2 ? shout_r : _out_xpr_length_T_10; // @[alu.scala 73:8]
  wire [31:0] _out_xpr_length_T_12 = io_fn == 4'hc | io_fn == 4'he ? {{31'd0}, less} : _out_xpr_length_T_11; // @[alu.scala 72:8]
  assign io_out = io_fn == 4'h0 | io_fn == 4'ha ? sum : _out_xpr_length_T_12; // @[alu.scala 71:8]
  assign io_adder_out = io_in1 + _sum_T_3; // @[alu.scala 50:20]
endmodule