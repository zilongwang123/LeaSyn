//`define _EXTERNALMEMORY_

module ibex_top (
	clk_i,
	rst_ni,
	test_en_i,
	ram_cfg_i,
	hart_id_i,
	boot_addr_i,
	`ifdef _EXTERNALMEMORY_
		instr_req_o,
		instr_gnt_i,
		instr_rvalid_i,
		instr_addr_o,
		instr_rdata_i,
		instr_rdata_intg_i,
		instr_err_i,
		data_req_o,
		data_gnt_i,
		data_rvalid_i,
		data_we_o,
		data_be_o,
		data_addr_o,
		data_wdata_o,
		data_wdata_intg_o,
		data_rdata_i,
		data_rdata_intg_i,
		data_err_i,
	`endif
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	irq_nm_i,
	scramble_key_valid_i,
	scramble_key_i,
	scramble_nonce_i,
	scramble_req_o,
	debug_req_i,
	crash_dump_o,
	double_fault_seen_o,
	rvfi_valid,
	rvfi_order,
	rvfi_insn,
	rvfi_trap,
	rvfi_halt,
	rvfi_intr,
	rvfi_mode,
	rvfi_ixl,
	rvfi_rs1_addr,
	rvfi_rs2_addr,
	rvfi_rs3_addr,
	rvfi_rs1_rdata,
	rvfi_rs2_rdata,
	rvfi_rs3_rdata,
	rvfi_rd_addr,
	rvfi_rd_wdata,
	rvfi_pc_rdata,
	rvfi_pc_wdata,
	rvfi_mem_addr,
	rvfi_mem_rmask,
	rvfi_mem_wmask,
	rvfi_mem_rdata,
	rvfi_mem_wdata,
	// rvfi_ext_mip,
	// rvfi_ext_nmi,
	// rvfi_ext_nmi_int,
	// rvfi_ext_debug_req,
	// rvfi_ext_debug_mode,
	// rvfi_ext_rf_wr_suppress,
	// rvfi_ext_mcycle,
	// rvfi_ext_mhpmcounters,
	// rvfi_ext_mhpmcountersh,
	// rvfi_ext_ic_scr_key_valid,
	fetch_enable_i,
	alert_minor_o,
	alert_major_internal_o,
	alert_major_bus_o,
	core_sleep_o,
	scan_rst_ni,
);
	parameter [0:0] PMPEnable = 1'b0;
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumRegions = 4;
	parameter [31:0] MHPMCounterNum = 0;
	parameter [31:0] MHPMCounterWidth = 40;
	parameter [0:0] RV32E = 1'b0;
	parameter integer RV32M = 32'sd2;
	parameter integer RV32B = 32'sd0;
	parameter integer RegFile = 32'sd0;
	parameter [0:0] BranchTargetALU = 1'b0;
	parameter [0:0] WritebackStage = 1'b0;
	parameter [0:0] ICache = 1'b0;
	parameter [0:0] ICacheECC = 1'b0;
	parameter [0:0] BranchPredictor = 1'b0;
	parameter [0:0] DbgTriggerEn = 1'b0;
	parameter [31:0] DbgHwBreakNum = 1;
	parameter [0:0] SecureIbex = 1'b0;
	parameter [0:0] ICacheScramble = 1'b0;
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	localparam [31:0] ibex_pkg_SCRAMBLE_KEY_W = 128;
	localparam [127:0] ibex_pkg_RndCnstIbexKeyDefault = 128'h14e8cecae3040d5e12286bb3cc113298;
	parameter [127:0] RndCnstIbexKey = ibex_pkg_RndCnstIbexKeyDefault;
	localparam [31:0] ibex_pkg_SCRAMBLE_NONCE_W = 64;
	localparam [63:0] ibex_pkg_RndCnstIbexNonceDefault = 64'hf79780bc735f3843;
	parameter [63:0] RndCnstIbexNonce = ibex_pkg_RndCnstIbexNonceDefault;
	input wire clk_i;
	input wire rst_ni;
	input wire test_en_i;
	input wire [9:0] ram_cfg_i;
	input wire [31:0] hart_id_i;
	input wire [31:0] boot_addr_i;
	`ifdef _EXTERNALMEMORY_
		output wire instr_req_o;
		input wire instr_gnt_i;
		input wire instr_rvalid_i;
		output wire [31:0] instr_addr_o;
		input wire [31:0] instr_rdata_i;
		input wire [6:0] instr_rdata_intg_i;
		input wire instr_err_i;
		output wire data_req_o;
		input wire data_gnt_i;
		input wire data_rvalid_i;
		output wire data_we_o;
		output wire [3:0] data_be_o;
		output wire [31:0] data_addr_o;
		output wire [31:0] data_wdata_o;
		output wire [6:0] data_wdata_intg_o;
		input wire [31:0] data_rdata_i;
		input wire [6:0] data_rdata_intg_i;
		input wire data_err_i;
	`else
		wire instr_req_o;
		wire instr_gnt_i;//
	 	wire instr_rvalid_i;//
		wire [31:0] instr_addr_o;
		wire [31:0] instr_rdata_i;
		wire [6:0] instr_rdata_intg_i = 0;// not used
		wire instr_err_i = 0;//
		wire data_req_o;
		wire data_gnt_i;//set to high if the writing is finished
		wire data_rvalid_i;// indicates that the read date and err signal are valid
		wire data_we_o;// high for writes, low for reads
		wire [3:0] data_be_o;//
		wire [31:0] data_addr_o;
		wire [31:0] data_wdata_o;
		wire [6:0] data_wdata_intg_o = 0;// not used
		wire [31:0] data_rdata_i;
		wire [6:0] data_rdata_intg_i = 0;// not used
		wire data_err_i = 0;//
		ibex_imem ibex_imem(
				.clk(clk_i),
				.sram_req(instr_req_o),
				.sram_gnt(instr_gnt_i),
				.sram_rvalid(instr_rvalid_i),
				.sram_addr(instr_addr_o[11:2]),
				.sram_rdata(instr_rdata_i),
				.pc_ctr(pc_ctr),
				.instr_ctr(instr_ctr),
				.rvfi_pc_ctr(rvfi_pc_ctr),
				.rvfi_instr_ctr(rvfi_instr_ctr),
				.pc_id(pc_id),
		);
		ibex_dmem ibex_dmem(
				.clk(clk_i),
				.sram_req(data_req_o),
				.sram_gnt(data_gnt_i),
				.sram_rvalid(data_rvalid_i),
				.sram_we(data_we_o),
				.sram_be(data_be_o),
				.sram_addr(data_addr_o[11:2]),
				.sram_wdata(data_wdata_o),
				.sram_rdata(data_rdata_i),
				.lsu_addr_ctr(lsu_addr_ctr),
		);
	`endif
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [14:0] irq_fast_i;
	input wire irq_nm_i;
	input wire scramble_key_valid_i;
	input wire [127:0] scramble_key_i;
	input wire [63:0] scramble_nonce_i;
	output wire scramble_req_o;
	input wire debug_req_i;
	output wire [159:0] crash_dump_o;
	output wire double_fault_seen_o;
	output wire rvfi_valid;
	output wire [63:0] rvfi_order;
	output wire [31:0] rvfi_insn;
	output wire rvfi_trap;
	output wire rvfi_halt;
	output wire rvfi_intr;
	output wire [1:0] rvfi_mode;
	output wire [1:0] rvfi_ixl;
	output wire [4:0] rvfi_rs1_addr;
	output wire [4:0] rvfi_rs2_addr;
	output wire [4:0] rvfi_rs3_addr;
	output wire [31:0] rvfi_rs1_rdata;
	output wire [31:0] rvfi_rs2_rdata;
	output wire [31:0] rvfi_rs3_rdata;
	output wire [4:0] rvfi_rd_addr;
	output wire [31:0] rvfi_rd_wdata;
	output wire [31:0] rvfi_pc_rdata;
	output wire [31:0] rvfi_pc_wdata;
	output wire [31:0] rvfi_mem_addr;
	output wire [3:0] rvfi_mem_rmask;
	output wire [3:0] rvfi_mem_wmask;
	output wire [31:0] rvfi_mem_rdata;
	output wire [31:0] rvfi_mem_wdata;
	// output wire [31:0] rvfi_ext_mip;
	// output wire rvfi_ext_nmi;
	// output wire rvfi_ext_nmi_int;
	// output wire rvfi_ext_debug_req;
	// output wire rvfi_ext_debug_mode;
	// output wire rvfi_ext_rf_wr_suppress;
	// output wire [63:0] rvfi_ext_mcycle;
	// output wire [319:0] rvfi_ext_mhpmcounters;
	// output wire [319:0] rvfi_ext_mhpmcountersh;
	// output wire rvfi_ext_ic_scr_key_valid;
	input wire [3:0] fetch_enable_i;
	output wire alert_minor_o;
	output wire alert_major_internal_o;
	output wire alert_major_bus_o;
	output wire core_sleep_o;
	input wire scan_rst_ni;
	localparam [0:0] Lockstep = SecureIbex;
	localparam [0:0] ResetAll = Lockstep;
	localparam [0:0] DummyInstructions = SecureIbex;
	localparam [0:0] RegFileECC = SecureIbex;
	localparam [0:0] RegFileWrenCheck = SecureIbex;
	localparam [31:0] RegFileDataWidth = (RegFileECC ? 39 : 32);
	localparam [0:0] MemECC = SecureIbex;
	localparam [31:0] MemDataWidth = (MemECC ? 39 : 32);
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	localparam [31:0] BusSizeECC = (ICacheECC ? 39 : ibex_pkg_BUS_SIZE);
	localparam [31:0] ibex_pkg_BUS_BYTES = 4;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_LINE_BEATS = ibex_pkg_IC_LINE_BYTES / ibex_pkg_BUS_BYTES;
	localparam [31:0] LineSizeECC = BusSizeECC * ibex_pkg_IC_LINE_BEATS;
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	localparam [31:0] TagSizeECC = (ICacheECC ? ibex_pkg_IC_TAG_SIZE + 6 : ibex_pkg_IC_TAG_SIZE);
	localparam [31:0] NumAddrScrRounds = (ICacheScramble ? 2 : 0);
	localparam [31:0] NumDiffRounds = NumAddrScrRounds;
	wire clk;
	wire [3:0] core_busy_d;
	reg [3:0] core_busy_q;
	wire clock_en;
	wire irq_pending;
	wire dummy_instr_id;
	wire dummy_instr_wb;
	wire [4:0] rf_raddr_a;
	wire [4:0] rf_raddr_b;
	wire [4:0] rf_waddr_wb;
	wire rf_we_wb;
	wire [RegFileDataWidth - 1:0] rf_wdata_wb_ecc;
	wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc;
	wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc_buf;
	wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc;
	wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc_buf;
	wire [MemDataWidth - 1:0] data_wdata_core;
	wire [MemDataWidth - 1:0] data_rdata_core;
	wire [MemDataWidth - 1:0] instr_rdata_core;
	wire [1:0] ic_tag_req;
	wire ic_tag_write;
	wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr;
	wire [TagSizeECC - 1:0] ic_tag_wdata;
	wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata;
	wire [1:0] ic_data_req;
	wire ic_data_write;
	wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr;
	wire [LineSizeECC - 1:0] ic_data_wdata;
	wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata;
	wire ic_scr_key_req;
	wire core_alert_major_internal;
	wire core_alert_major_bus;
	wire core_alert_minor;
	wire lockstep_alert_major_internal;
	wire lockstep_alert_major_bus;
	wire lockstep_alert_minor;
	reg [127:0] scramble_key_q;
	reg [63:0] scramble_nonce_q;
	wire scramble_key_valid_d;
	reg scramble_key_valid_q;
	wire scramble_req_d;
	reg scramble_req_q;
	wire [3:0] fetch_enable_buf;
	localparam [3:0] ibex_pkg_IbexMuBiOff = 4'b1010;
	// generate
	// 	if (SecureIbex) begin : g_clock_en_secure
	// 		prim_generic_flop #(
	// 			.Width(4),
	// 			.ResetValue(ibex_pkg_IbexMuBiOff)
	// 		) u_prim_core_busy_flop(
	// 			.clk_i(clk_i),
	// 			.rst_ni(rst_ni),
	// 			.d_i(core_busy_d),
	// 			.q_o(core_busy_q)
	// 		);
	// 		assign clock_en = (((core_busy_q != ibex_pkg_IbexMuBiOff) | debug_req_i) | irq_pending) | irq_nm_i;
	// 	end
	// 	else begin : g_clock_en_non_secure
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					core_busy_q <= ibex_pkg_IbexMuBiOff;
				else
					core_busy_q <= core_busy_d;
			assign clock_en = ((core_busy_q[0] | debug_req_i) | irq_pending) | irq_nm_i;
			wire unused_core_busy;
			assign unused_core_busy = ^core_busy_q[3:1];
	// 	end
	// endgenerate
	assign core_sleep_o = ~clock_en;
	prim_clock_gating prim_clock_gating(
		.clk_i(clk_i),
		.en_i(clock_en),
		.test_en_i(test_en_i),
		.clk_o(clk)
	);
	prim_generic_buf #(.Width(4)) u_fetch_enable_buf(
		.in_i(fetch_enable_i),
		.out_o(fetch_enable_buf)
	);
	prim_generic_buf #(.Width(RegFileDataWidth)) u_rf_rdata_a_ecc_buf(
		.in_i(rf_rdata_a_ecc),
		.out_o(rf_rdata_a_ecc_buf)
	);
	prim_generic_buf #(.Width(RegFileDataWidth)) u_rf_rdata_b_ecc_buf(
		.in_i(rf_rdata_b_ecc),
		.out_o(rf_rdata_b_ecc_buf)
	);
	assign data_rdata_core[31:0] = data_rdata_i;
	assign instr_rdata_core[31:0] = instr_rdata_i;
	// generate
	// 	if (MemECC) begin : gen_mem_rdata_ecc
	// 		assign data_rdata_core[38:32] = data_rdata_intg_i;
	// 		assign instr_rdata_core[38:32] = instr_rdata_intg_i;
	// 	end
	// 	else begin : gen_non_mem_rdata_ecc
			wire unused_intg;
			assign unused_intg = ^{instr_rdata_intg_i, data_rdata_intg_i};
	// 	end
	// endgenerate
	ibex_core #(
		.PMPEnable(PMPEnable),
		.PMPGranularity(PMPGranularity),
		.PMPNumRegions(PMPNumRegions),
		.MHPMCounterNum(MHPMCounterNum),
		.MHPMCounterWidth(MHPMCounterWidth),
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU),
		.ICache(ICache),
		.ICacheECC(ICacheECC),
		.BusSizeECC(BusSizeECC),
		.TagSizeECC(TagSizeECC),
		.LineSizeECC(LineSizeECC),
		.BranchPredictor(BranchPredictor),
		.DbgTriggerEn(DbgTriggerEn),
		.DbgHwBreakNum(DbgHwBreakNum),
		.WritebackStage(WritebackStage),
		.ResetAll(ResetAll),
		.RndCnstLfsrSeed(RndCnstLfsrSeed),
		.RndCnstLfsrPerm(RndCnstLfsrPerm),
		.SecureIbex(SecureIbex),
		.DummyInstructions(DummyInstructions),
		.RegFileECC(RegFileECC),
		.RegFileDataWidth(RegFileDataWidth),
		.MemECC(MemECC),
		.MemDataWidth(MemDataWidth),
		.DmHaltAddr(DmHaltAddr),
		.DmExceptionAddr(DmExceptionAddr)
	) ibex_core(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.hart_id_i(hart_id_i),
		.boot_addr_i(boot_addr_i),
		.instr_req_o(instr_req_o),
		.instr_gnt_i(instr_gnt_i),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_addr_o(instr_addr_o),
		.instr_rdata_i(instr_rdata_core),
		.instr_err_i(instr_err_i),
		.data_req_o(data_req_o),
		.data_gnt_i(data_gnt_i),
		.data_rvalid_i(data_rvalid_i),
		.data_we_o(data_we_o),
		.data_be_o(data_be_o),
		.data_addr_o(data_addr_o),
		.data_wdata_o(data_wdata_core),
		.data_rdata_i(data_rdata_core),
		.data_err_i(data_err_i),
		.dummy_instr_id_o(dummy_instr_id),
		.dummy_instr_wb_o(dummy_instr_wb),
		.rf_raddr_a_o(rf_raddr_a),
		.rf_raddr_b_o(rf_raddr_b),
		.rf_waddr_wb_o(rf_waddr_wb),
		.rf_we_wb_o(rf_we_wb),
		.rf_wdata_wb_ecc_o(rf_wdata_wb_ecc),
		.rf_rdata_a_ecc_i(rf_rdata_a_ecc_buf),
		.rf_rdata_b_ecc_i(rf_rdata_b_ecc_buf),
		.ic_tag_req_o(ic_tag_req),
		.ic_tag_write_o(ic_tag_write),
		.ic_tag_addr_o(ic_tag_addr),
		.ic_tag_wdata_o(ic_tag_wdata),
		.ic_tag_rdata_i(ic_tag_rdata),
		.ic_data_req_o(ic_data_req),
		.ic_data_write_o(ic_data_write),
		.ic_data_addr_o(ic_data_addr),
		.ic_data_wdata_o(ic_data_wdata),
		.ic_data_rdata_i(ic_data_rdata),
		.ic_scr_key_valid_i(scramble_key_valid_q),
		.ic_scr_key_req_o(ic_scr_key_req),
		.irq_software_i(irq_software_i),
		.irq_timer_i(irq_timer_i),
		.irq_external_i(irq_external_i),
		.irq_fast_i(irq_fast_i),
		.irq_nm_i(irq_nm_i),
		.irq_pending_o(irq_pending),
		.debug_req_i(debug_req_i),
		.crash_dump_o(crash_dump_o),
		.double_fault_seen_o(double_fault_seen_o),
		.rvfi_valid(rvfi_valid),
		.rvfi_order(rvfi_order),
		.rvfi_insn(rvfi_insn),
		.rvfi_trap(rvfi_trap),
		.rvfi_halt(rvfi_halt),
		.rvfi_intr(rvfi_intr),
		.rvfi_mode(rvfi_mode),
		.rvfi_ixl(rvfi_ixl),
		.rvfi_rs1_addr(rvfi_rs1_addr),
		.rvfi_rs2_addr(rvfi_rs2_addr),
		.rvfi_rs3_addr(rvfi_rs3_addr),
		.rvfi_rs1_rdata(rvfi_rs1_rdata),
		.rvfi_rs2_rdata(rvfi_rs2_rdata),
		.rvfi_rs3_rdata(rvfi_rs3_rdata),
		.rvfi_rd_addr(rvfi_rd_addr),
		.rvfi_rd_wdata(rvfi_rd_wdata),
		.rvfi_pc_rdata(rvfi_pc_rdata),
		.rvfi_pc_wdata(rvfi_pc_wdata),
		.rvfi_mem_addr(rvfi_mem_addr),
		.rvfi_mem_rmask(rvfi_mem_rmask),
		.rvfi_mem_wmask(rvfi_mem_wmask),
		.rvfi_mem_rdata(rvfi_mem_rdata),
		.rvfi_mem_wdata(rvfi_mem_wdata),
		// .rvfi_ext_mip(rvfi_ext_mip),
		// .rvfi_ext_nmi(rvfi_ext_nmi),
		// .rvfi_ext_nmi_int(rvfi_ext_nmi_int),
		// .rvfi_ext_debug_req(rvfi_ext_debug_req),
		// .rvfi_ext_debug_mode(rvfi_ext_debug_mode),
		// .rvfi_ext_rf_wr_suppress(rvfi_ext_rf_wr_suppress),
		// .rvfi_ext_mcycle(rvfi_ext_mcycle),
		// .rvfi_ext_mhpmcounters(rvfi_ext_mhpmcounters),
		// .rvfi_ext_mhpmcountersh(rvfi_ext_mhpmcountersh),
		// .rvfi_ext_ic_scr_key_valid(rvfi_ext_ic_scr_key_valid),
		.fetch_enable_i(fetch_enable_buf),
		.alert_minor_o(core_alert_minor),
		.alert_major_internal_o(core_alert_major_internal),
		.alert_major_bus_o(core_alert_major_bus),
		.core_busy_o(core_busy_d),
		//// for contract
		.pc_ctr(pc_ctr),
		.instr_ctr(instr_ctr),
		.rvfi_pc_ctr(rvfi_pc_ctr),
		.rvfi_instr_ctr(rvfi_instr_ctr),
		.pc_id(pc_id),
		.rf_raddr_a_o_ctr(rf_raddr_a_o_ctr),
		.rf_raddr_b_o_ctr(rf_raddr_b_o_ctr),
		.rf_raddr_b_o_ctr_id(rf_raddr_b_o_ctr_id),
		.rf_raddr_a_o_ctr_id(rf_raddr_a_o_ctr_id),
		.rf_rdata_a_fwd_ctr(rf_rdata_a_fwd_ctr),
		.rf_rdata_b_fwd_ctr(rf_rdata_b_fwd_ctr),
		.rf_rdata_b_fwd_ctr_id(rf_rdata_b_fwd_ctr_id),
		.rf_rdata_a_fwd_ctr_id(rf_rdata_a_fwd_ctr_id),
		.lsu_addr_ctr(lsu_addr_ctr),
	);
	//// for contract
	wire [31:0] pc_ctr;
	wire [31:0] instr_ctr;
	wire [31:0] rvfi_pc_ctr;
	wire [31:0] rvfi_instr_ctr;
	wire [31:0] pc_id;
	wire [4:0]  rf_raddr_a_o_ctr;
	wire [4:0]  rf_raddr_b_o_ctr;
	wire [4:0]  rf_raddr_b_o_ctr_id;
	wire [4:0]  rf_raddr_a_o_ctr_id;
	wire [31:0]	rf_rdata_a_fwd_ctr;
	wire [31:0]	rf_rdata_b_fwd_ctr;
	wire [31:0]	rf_rdata_b_fwd_ctr_id;
	wire [31:0]	rf_rdata_a_fwd_ctr_id;
	wire [31:0] lsu_addr_ctr;




	wire rf_alert_major_internal;
	localparam [38:0] prim_secded_pkg_SecdedInv3932ZeroWord = 39'h2a00000000;
	function automatic [RegFileDataWidth - 1:0] sv2v_cast_E67BC;
		input reg [RegFileDataWidth - 1:0] inp;
		sv2v_cast_E67BC = inp;
	endfunction
	// generate
	// 	if (RegFile == 32'sd0) begin : gen_regfile_ff
			ibex_register_file_ff #(
				.RV32E(RV32E),
				.DataWidth(RegFileDataWidth),
				.DummyInstructions(DummyInstructions),
				.WrenCheck(RegFileWrenCheck),
				.WordZeroVal(sv2v_cast_E67BC(prim_secded_pkg_SecdedInv3932ZeroWord))
			) ibex_register_file_ff(
				.clk_i(clk),
				.rst_ni(rst_ni),
				.test_en_i(test_en_i),
				.dummy_instr_id_i(dummy_instr_id),
				.dummy_instr_wb_i(dummy_instr_wb),
				.raddr_a_i(rf_raddr_a),
				.rdata_a_o(rf_rdata_a_ecc),
				.raddr_b_i(rf_raddr_b),
				.rdata_b_o(rf_rdata_b_ecc),
				.waddr_a_i(rf_waddr_wb),
				.wdata_a_i(rf_wdata_wb_ecc),
				.we_a_i(rf_we_wb),
				.err_o(rf_alert_major_internal),
				.rf_raddr_a_o_ctr(rf_raddr_a_o_ctr),
				.rf_raddr_b_o_ctr(rf_raddr_b_o_ctr),
				.rf_raddr_b_o_ctr_id(rf_raddr_b_o_ctr_id),
				.rf_raddr_a_o_ctr_id(rf_raddr_a_o_ctr_id),
				.rf_rdata_a_fwd_ctr(rf_rdata_a_fwd_ctr),
				.rf_rdata_b_fwd_ctr(rf_rdata_b_fwd_ctr),
				.rf_rdata_b_fwd_ctr_id(rf_rdata_b_fwd_ctr_id),
				.rf_rdata_a_fwd_ctr_id(rf_rdata_a_fwd_ctr_id),
			);
		// end
		// else if (RegFile == 32'sd1) begin : gen_regfile_fpga
		// 	ibex_register_file_fpga #(
		// 		.RV32E(RV32E),
		// 		.DataWidth(RegFileDataWidth),
		// 		.DummyInstructions(DummyInstructions),
		// 		.WrenCheck(RegFileWrenCheck),
		// 		.WordZeroVal(sv2v_cast_E67BC(prim_secded_pkg_SecdedInv3932ZeroWord))
		// 	) ibex_register_file_fpga(
		// 		.clk_i(clk),
		// 		.rst_ni(rst_ni),
		// 		.test_en_i(test_en_i),
		// 		.dummy_instr_id_i(dummy_instr_id),
		// 		.dummy_instr_wb_i(dummy_instr_wb),
		// 		.raddr_a_i(rf_raddr_a),
		// 		.rdata_a_o(rf_rdata_a_ecc),
		// 		.raddr_b_i(rf_raddr_b),
		// 		.rdata_b_o(rf_rdata_b_ecc),
		// 		.waddr_a_i(rf_waddr_wb),
		// 		.wdata_a_i(rf_wdata_wb_ecc),
		// 		.we_a_i(rf_we_wb),
		// 		.err_o(rf_alert_major_internal)
		// 	);
		// end
		// else if (RegFile == 32'sd2) begin : gen_regfile_latch
		// 	ibex_register_file_latch #(
		// 		.RV32E(RV32E),
		// 		.DataWidth(RegFileDataWidth),
		// 		.DummyInstructions(DummyInstructions),
		// 		.WrenCheck(RegFileWrenCheck),
		// 		.WordZeroVal(sv2v_cast_E67BC(prim_secded_pkg_SecdedInv3932ZeroWord))
		// 	) ibex_register_file_latch(
		// 		.clk_i(clk),
		// 		.rst_ni(rst_ni),
		// 		.test_en_i(test_en_i),
		// 		.dummy_instr_id_i(dummy_instr_id),
		// 		.dummy_instr_wb_i(dummy_instr_wb),
		// 		.raddr_a_i(rf_raddr_a),
		// 		.rdata_a_o(rf_rdata_a_ecc),
		// 		.raddr_b_i(rf_raddr_b),
		// 		.rdata_b_o(rf_rdata_b_ecc),
		// 		.waddr_a_i(rf_waddr_wb),
		// 		.wdata_a_i(rf_wdata_wb_ecc),
		// 		.we_a_i(rf_we_wb),
		// 		.err_o(rf_alert_major_internal)
		// 	);
		// end
		// if (ICacheScramble) begin : gen_scramble
		// 	assign scramble_key_valid_d = (scramble_req_q ? scramble_key_valid_i : (ic_scr_key_req ? 1'b0 : scramble_key_valid_q));
		// 	always @(posedge clk_i or negedge rst_ni)
		// 		if (!rst_ni) begin
		// 			scramble_key_q <= RndCnstIbexKey;
		// 			scramble_nonce_q <= RndCnstIbexNonce;
		// 		end
		// 		else if (scramble_key_valid_i) begin
		// 			scramble_key_q <= scramble_key_i;
		// 			scramble_nonce_q <= scramble_nonce_i;
		// 		end
		// 	always @(posedge clk_i or negedge rst_ni)
		// 		if (!rst_ni) begin
		// 			scramble_key_valid_q <= 1'b1;
		// 			scramble_req_q <= 1'sb0;
		// 		end
		// 		else begin
		// 			scramble_key_valid_q <= scramble_key_valid_d;
		// 			scramble_req_q <= scramble_req_d;
		// 		end
		// 	assign scramble_req_d = (scramble_req_q ? ~scramble_key_valid_i : ic_scr_key_req);
		// 	assign scramble_req_o = scramble_req_q;
		// end
		// else begin : gen_noscramble
			reg unused_scramble_inputs = (((((((scramble_key_valid_i & |scramble_key_i) & |RndCnstIbexKey) & |scramble_nonce_i) & |RndCnstIbexNonce) & scramble_req_q) & ic_scr_key_req) & scramble_key_valid_d) & scramble_req_d;
			assign scramble_req_d = 1'b0;
			wire [1:1] sv2v_tmp_AE3A4;
			assign sv2v_tmp_AE3A4 = 1'b0;
			always @(*) scramble_req_q = sv2v_tmp_AE3A4;
			assign scramble_req_o = 1'b0;
			wire [128:1] sv2v_tmp_A2325;
			assign sv2v_tmp_A2325 = 1'sb0;
			always @(*) scramble_key_q = sv2v_tmp_A2325;
			wire [64:1] sv2v_tmp_70913;
			assign sv2v_tmp_70913 = 1'sb0;
			always @(*) scramble_nonce_q = sv2v_tmp_70913;
			wire [1:1] sv2v_tmp_92821;
			assign sv2v_tmp_92821 = 1'b1;
			always @(*) scramble_key_valid_q = sv2v_tmp_92821;
			assign scramble_key_valid_d = 1'b1;
	// 	end
	// endgenerate
	function automatic [TagSizeECC - 1:0] sv2v_cast_BD0FC;
		input reg [TagSizeECC - 1:0] inp;
		sv2v_cast_BD0FC = inp;
	endfunction
	function automatic [LineSizeECC - 1:0] sv2v_cast_F09E7;
		input reg [LineSizeECC - 1:0] inp;
		sv2v_cast_F09E7 = inp;
	endfunction
	// generate
	// 	if (ICache) begin : gen_rams
	// 		genvar way;
	// 		for (way = 0; way < ibex_pkg_IC_NUM_WAYS; way = way + 1) begin : gen_rams_inner
	// 			if (ICacheScramble) begin : gen_scramble_rams
	// 				prim_ram_1p_scr #(
	// 					.Width(TagSizeECC),
	// 					.Depth(ibex_pkg_IC_NUM_LINES),
	// 					.DataBitsPerMask(TagSizeECC),
	// 					.EnableParity(0),
	// 					.DiffWidth(TagSizeECC),
	// 					.NumAddrScrRounds(NumAddrScrRounds),
	// 					.NumDiffRounds(NumDiffRounds)
	// 				) tag_bank(
	// 					.clk_i(clk_i),
	// 					.rst_ni(rst_ni),
	// 					.key_valid_i(scramble_key_valid_q),
	// 					.key_i(scramble_key_q),
	// 					.nonce_i(scramble_nonce_q),
	// 					.req_i(ic_tag_req[way]),
	// 					.gnt_o(),
	// 					.write_i(ic_tag_write),
	// 					.addr_i(ic_tag_addr),
	// 					.wdata_i(ic_tag_wdata),
	// 					.wmask_i({TagSizeECC {1'b1}}),
	// 					.intg_error_i(1'b0),
	// 					.rdata_o(ic_tag_rdata[(1 - way) * TagSizeECC+:TagSizeECC]),
	// 					.rvalid_o(),
	// 					.raddr_o(),
	// 					.rerror_o(),
	// 					.cfg_i(ram_cfg_i)
	// 				);
	// 				prim_ram_1p_scr #(
	// 					.Width(LineSizeECC),
	// 					.Depth(ibex_pkg_IC_NUM_LINES),
	// 					.DataBitsPerMask(LineSizeECC),
	// 					.ReplicateKeyStream(1),
	// 					.EnableParity(0),
	// 					.DiffWidth(LineSizeECC),
	// 					.NumAddrScrRounds(NumAddrScrRounds),
	// 					.NumDiffRounds(NumDiffRounds)
	// 				) data_bank(
	// 					.clk_i(clk_i),
	// 					.rst_ni(rst_ni),
	// 					.key_valid_i(scramble_key_valid_q),
	// 					.key_i(scramble_key_q),
	// 					.nonce_i(scramble_nonce_q),
	// 					.req_i(ic_data_req[way]),
	// 					.gnt_o(),
	// 					.write_i(ic_data_write),
	// 					.addr_i(ic_data_addr),
	// 					.wdata_i(ic_data_wdata),
	// 					.wmask_i({LineSizeECC {1'b1}}),
	// 					.intg_error_i(1'b0),
	// 					.rdata_o(ic_data_rdata[(1 - way) * LineSizeECC+:LineSizeECC]),
	// 					.rvalid_o(),
	// 					.raddr_o(),
	// 					.rerror_o(),
	// 					.cfg_i(ram_cfg_i)
	// 				);
	// 			end
	// 			else begin : gen_noscramble_rams
	// 				prim_ram_1p #(
	// 					.Width(TagSizeECC),
	// 					.Depth(ibex_pkg_IC_NUM_LINES),
	// 					.DataBitsPerMask(TagSizeECC)
	// 				) tag_bank(
	// 					.clk_i(clk_i),
	// 					.req_i(ic_tag_req[way]),
	// 					.write_i(ic_tag_write),
	// 					.addr_i(ic_tag_addr),
	// 					.wdata_i(ic_tag_wdata),
	// 					.wmask_i({TagSizeECC {1'b1}}),
	// 					.rdata_o(ic_tag_rdata[(1 - way) * TagSizeECC+:TagSizeECC]),
	// 					.cfg_i(ram_cfg_i)
	// 				);
	// 				prim_ram_1p #(
	// 					.Width(LineSizeECC),
	// 					.Depth(ibex_pkg_IC_NUM_LINES),
	// 					.DataBitsPerMask(LineSizeECC)
	// 				) data_bank(
	// 					.clk_i(clk_i),
	// 					.req_i(ic_data_req[way]),
	// 					.write_i(ic_data_write),
	// 					.addr_i(ic_data_addr),
	// 					.wdata_i(ic_data_wdata),
	// 					.wmask_i({LineSizeECC {1'b1}}),
	// 					.rdata_o(ic_data_rdata[(1 - way) * LineSizeECC+:LineSizeECC]),
	// 					.cfg_i(ram_cfg_i)
	// 				);
	// 			end
	// 		end
	// 	end
	// 	else begin : gen_norams
			wire [9:0] unused_ram_cfg;
			wire unused_ram_inputs;
			assign unused_ram_cfg = ram_cfg_i;
			assign unused_ram_inputs = ((((((((((((|ic_tag_req & ic_tag_write) & |ic_tag_addr) & |ic_tag_wdata) & |ic_data_req) & ic_data_write) & |ic_data_addr) & |ic_data_wdata) & |scramble_key_q) & |scramble_nonce_q) & scramble_key_valid_q) & scramble_key_valid_d) & |scramble_nonce_q) & |NumAddrScrRounds;
			assign ic_tag_rdata = {ibex_pkg_IC_NUM_WAYS {sv2v_cast_BD0FC('b0)}};
			assign ic_data_rdata = {ibex_pkg_IC_NUM_WAYS {sv2v_cast_F09E7('b0)}};
	// 	end
	// endgenerate
	assign data_wdata_o = data_wdata_core[31:0];
	// generate
	// 	if (MemECC) begin : gen_mem_wdata_ecc
	// 		prim_generic_buf #(.Width(7)) u_prim_generic_buf_data_wdata_intg(
	// 			.in_i(data_wdata_core[38:32]),
	// 			.out_o(data_wdata_intg_o)
	// 		);
	// 	end
	// 	else begin : gen_no_mem_ecc
			assign data_wdata_intg_o = 1'sb0;
		// end
		// if (Lockstep) begin : gen_lockstep
		// 	localparam signed [31:0] NumBufferBits = ((((((((((((((((99 + MemDataWidth) + 41) + MemDataWidth) + MemDataWidth) + 19) + RegFileDataWidth) + RegFileDataWidth) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 192;
		// 	wire [NumBufferBits - 1:0] buf_in;
		// 	wire [NumBufferBits - 1:0] buf_out;
		// 	wire [31:0] hart_id_local;
		// 	wire [31:0] boot_addr_local;
		// 	wire instr_req_local;
		// 	wire instr_gnt_local;
		// 	wire instr_rvalid_local;
		// 	wire [31:0] instr_addr_local;
		// 	wire [MemDataWidth - 1:0] instr_rdata_local;
		// 	wire instr_err_local;
		// 	wire data_req_local;
		// 	wire data_gnt_local;
		// 	wire data_rvalid_local;
		// 	wire data_we_local;
		// 	wire [3:0] data_be_local;
		// 	wire [31:0] data_addr_local;
		// 	wire [MemDataWidth - 1:0] data_wdata_local;
		// 	wire [MemDataWidth - 1:0] data_rdata_local;
		// 	wire data_err_local;
		// 	wire dummy_instr_id_local;
		// 	wire dummy_instr_wb_local;
		// 	wire [4:0] rf_raddr_a_local;
		// 	wire [4:0] rf_raddr_b_local;
		// 	wire [4:0] rf_waddr_wb_local;
		// 	wire rf_we_wb_local;
		// 	wire [RegFileDataWidth - 1:0] rf_wdata_wb_ecc_local;
		// 	wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc_local;
		// 	wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc_local;
		// 	wire [1:0] ic_tag_req_local;
		// 	wire ic_tag_write_local;
		// 	wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_local;
		// 	wire [TagSizeECC - 1:0] ic_tag_wdata_local;
		// 	wire [1:0] ic_data_req_local;
		// 	wire ic_data_write_local;
		// 	wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_local;
		// 	wire [LineSizeECC - 1:0] ic_data_wdata_local;
		// 	wire scramble_key_valid_local;
		// 	wire ic_scr_key_req_local;
		// 	wire irq_software_local;
		// 	wire irq_timer_local;
		// 	wire irq_external_local;
		// 	wire [14:0] irq_fast_local;
		// 	wire irq_nm_local;
		// 	wire irq_pending_local;
		// 	wire debug_req_local;
		// 	wire [159:0] crash_dump_local;
		// 	wire double_fault_seen_local;
		// 	wire [3:0] fetch_enable_local;
		// 	wire [3:0] core_busy_local;
		// 	assign buf_in = {hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_core, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_core, data_rdata_core, data_err_i, dummy_instr_id, dummy_instr_wb, rf_raddr_a, rf_raddr_b, rf_waddr_wb, rf_we_wb, rf_wdata_wb_ecc, rf_rdata_a_ecc, rf_rdata_b_ecc, ic_tag_req, ic_tag_write, ic_tag_addr, ic_tag_wdata, ic_data_req, ic_data_write, ic_data_addr, ic_data_wdata, scramble_key_valid_q, ic_scr_key_req, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, irq_nm_i, irq_pending, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, core_busy_d};
		// 	assign {hart_id_local, boot_addr_local, instr_req_local, instr_gnt_local, instr_rvalid_local, instr_addr_local, instr_rdata_local, instr_err_local, data_req_local, data_gnt_local, data_rvalid_local, data_we_local, data_be_local, data_addr_local, data_wdata_local, data_rdata_local, data_err_local, dummy_instr_id_local, dummy_instr_wb_local, rf_raddr_a_local, rf_raddr_b_local, rf_waddr_wb_local, rf_we_wb_local, rf_wdata_wb_ecc_local, rf_rdata_a_ecc_local, rf_rdata_b_ecc_local, ic_tag_req_local, ic_tag_write_local, ic_tag_addr_local, ic_tag_wdata_local, ic_data_req_local, ic_data_write_local, ic_data_addr_local, ic_data_wdata_local, scramble_key_valid_local, ic_scr_key_req_local, irq_software_local, irq_timer_local, irq_external_local, irq_fast_local, irq_nm_local, irq_pending_local, debug_req_local, crash_dump_local, double_fault_seen_local, fetch_enable_local, core_busy_local} = buf_out;
		// 	prim_generic_buf #(.Width(NumBufferBits)) u_signals_prim_generic_buf(
		// 		.in_i(buf_in),
		// 		.out_o(buf_out)
		// 	);
		// 	wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_local;
		// 	wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_local;
		// 	genvar k;
		// 	for (k = 0; k < ibex_pkg_IC_NUM_WAYS; k = k + 1) begin : gen_ways
		// 		prim_generic_buf #(.Width(TagSizeECC)) u_tag_prim_generic_buf(
		// 			.in_i(ic_tag_rdata[(1 - k) * TagSizeECC+:TagSizeECC]),
		// 			.out_o(ic_tag_rdata_local[(1 - k) * TagSizeECC+:TagSizeECC])
		// 		);
		// 		prim_generic_buf #(.Width(LineSizeECC)) u_data_prim_generic_buf(
		// 			.in_i(ic_data_rdata[(1 - k) * LineSizeECC+:LineSizeECC]),
		// 			.out_o(ic_data_rdata_local[(1 - k) * LineSizeECC+:LineSizeECC])
		// 		);
		// 	end
		// 	wire lockstep_alert_minor_local;
		// 	wire lockstep_alert_major_internal_local;
		// 	wire lockstep_alert_major_bus_local;
		// 	ibex_lockstep #(
		// 		.PMPEnable(PMPEnable),
		// 		.PMPGranularity(PMPGranularity),
		// 		.PMPNumRegions(PMPNumRegions),
		// 		.MHPMCounterNum(MHPMCounterNum),
		// 		.MHPMCounterWidth(MHPMCounterWidth),
		// 		.RV32E(RV32E),
		// 		.RV32M(RV32M),
		// 		.RV32B(RV32B),
		// 		.BranchTargetALU(BranchTargetALU),
		// 		.ICache(ICache),
		// 		.ICacheECC(ICacheECC),
		// 		.BusSizeECC(BusSizeECC),
		// 		.TagSizeECC(TagSizeECC),
		// 		.LineSizeECC(LineSizeECC),
		// 		.BranchPredictor(BranchPredictor),
		// 		.DbgTriggerEn(DbgTriggerEn),
		// 		.DbgHwBreakNum(DbgHwBreakNum),
		// 		.WritebackStage(WritebackStage),
		// 		.ResetAll(ResetAll),
		// 		.RndCnstLfsrSeed(RndCnstLfsrSeed),
		// 		.RndCnstLfsrPerm(RndCnstLfsrPerm),
		// 		.SecureIbex(SecureIbex),
		// 		.DummyInstructions(DummyInstructions),
		// 		.RegFileECC(RegFileECC),
		// 		.RegFileDataWidth(RegFileDataWidth),
		// 		.MemECC(MemECC),
		// 		.DmHaltAddr(DmHaltAddr),
		// 		.DmExceptionAddr(DmExceptionAddr)
		// 	) u_ibex_lockstep(
		// 		.clk_i(clk),
		// 		.rst_ni(rst_ni),
		// 		.hart_id_i(hart_id_local),
		// 		.boot_addr_i(boot_addr_local),
		// 		.instr_req_i(instr_req_local),
		// 		.instr_gnt_i(instr_gnt_local),
		// 		.instr_rvalid_i(instr_rvalid_local),
		// 		.instr_addr_i(instr_addr_local),
		// 		.instr_rdata_i(instr_rdata_local),
		// 		.instr_err_i(instr_err_local),
		// 		.data_req_i(data_req_local),
		// 		.data_gnt_i(data_gnt_local),
		// 		.data_rvalid_i(data_rvalid_local),
		// 		.data_we_i(data_we_local),
		// 		.data_be_i(data_be_local),
		// 		.data_addr_i(data_addr_local),
		// 		.data_wdata_i(data_wdata_local),
		// 		.data_rdata_i(data_rdata_local),
		// 		.data_err_i(data_err_local),
		// 		.dummy_instr_id_i(dummy_instr_id_local),
		// 		.dummy_instr_wb_i(dummy_instr_wb_local),
		// 		.rf_raddr_a_i(rf_raddr_a_local),
		// 		.rf_raddr_b_i(rf_raddr_b_local),
		// 		.rf_waddr_wb_i(rf_waddr_wb_local),
		// 		.rf_we_wb_i(rf_we_wb_local),
		// 		.rf_wdata_wb_ecc_i(rf_wdata_wb_ecc_local),
		// 		.rf_rdata_a_ecc_i(rf_rdata_a_ecc_local),
		// 		.rf_rdata_b_ecc_i(rf_rdata_b_ecc_local),
		// 		.ic_tag_req_i(ic_tag_req_local),
		// 		.ic_tag_write_i(ic_tag_write_local),
		// 		.ic_tag_addr_i(ic_tag_addr_local),
		// 		.ic_tag_wdata_i(ic_tag_wdata_local),
		// 		.ic_tag_rdata_i(ic_tag_rdata_local),
		// 		.ic_data_req_i(ic_data_req_local),
		// 		.ic_data_write_i(ic_data_write_local),
		// 		.ic_data_addr_i(ic_data_addr_local),
		// 		.ic_data_wdata_i(ic_data_wdata_local),
		// 		.ic_data_rdata_i(ic_data_rdata_local),
		// 		.ic_scr_key_valid_i(scramble_key_valid_local),
		// 		.ic_scr_key_req_i(ic_scr_key_req_local),
		// 		.irq_software_i(irq_software_local),
		// 		.irq_timer_i(irq_timer_local),
		// 		.irq_external_i(irq_external_local),
		// 		.irq_fast_i(irq_fast_local),
		// 		.irq_nm_i(irq_nm_local),
		// 		.irq_pending_i(irq_pending_local),
		// 		.debug_req_i(debug_req_local),
		// 		.crash_dump_i(crash_dump_local),
		// 		.double_fault_seen_i(double_fault_seen_local),
		// 		.fetch_enable_i(fetch_enable_local),
		// 		.alert_minor_o(lockstep_alert_minor_local),
		// 		.alert_major_internal_o(lockstep_alert_major_internal_local),
		// 		.alert_major_bus_o(lockstep_alert_major_bus_local),
		// 		.core_busy_i(core_busy_local),
		// 		.test_en_i(test_en_i),
		// 		.scan_rst_ni(scan_rst_ni)
		// 	);
		// 	prim_generic_buf u_prim_generic_buf_alert_minor(
		// 		.in_i(lockstep_alert_minor_local),
		// 		.out_o(lockstep_alert_minor)
		// 	);
		// 	prim_generic_buf u_prim_generic_buf_alert_major_internal(
		// 		.in_i(lockstep_alert_major_internal_local),
		// 		.out_o(lockstep_alert_major_internal)
		// 	);
		// 	prim_generic_buf u_prim_generic_buf_alert_major_bus(
		// 		.in_i(lockstep_alert_major_bus_local),
		// 		.out_o(lockstep_alert_major_bus)
		// 	);
		// end
		// else begin : gen_no_lockstep
			assign lockstep_alert_major_internal = 1'b0;
			assign lockstep_alert_major_bus = 1'b0;
			assign lockstep_alert_minor = 1'b0;
			wire unused_scan;
			assign unused_scan = scan_rst_ni;
	// 	end
	// endgenerate
	assign alert_major_internal_o = (core_alert_major_internal | lockstep_alert_major_internal) | rf_alert_major_internal;
	assign alert_major_bus_o = core_alert_major_bus | lockstep_alert_major_bus;
	assign alert_minor_o = core_alert_minor | lockstep_alert_minor;
endmodule
